//CAvium CA module testbench